//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.05
//Part Number: GW1NSR-LV4CQN48PC7/I6
//Device: GW1NSR-4C
//Created Time: Thu Feb 09 12:27:17 2023

module Gowin_ROM (dout, clk, oce, ce, reset, wre, ad);

output [11:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [9:0] ad;

wire [19:0] rom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

ROM rom_inst_0 (
    .DO({rom_inst_0_dout_w[19:0],dout[11:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam rom_inst_0.READ_MODE = 1'b0;
defparam rom_inst_0.BIT_WIDTH = 16;
defparam rom_inst_0.BLK_SEL = 3'b000;
defparam rom_inst_0.RESET_MODE = "ASYNC";
defparam rom_inst_0.INIT_RAM_00 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
defparam rom_inst_0.INIT_RAM_01 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
defparam rom_inst_0.INIT_RAM_02 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
defparam rom_inst_0.INIT_RAM_03 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
defparam rom_inst_0.INIT_RAM_04 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
defparam rom_inst_0.INIT_RAM_05 = 256'h000000000000000000000F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
defparam rom_inst_0.INIT_RAM_06 = 256'h000000000000000000000F0F0F0F0F0F0F0F0000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_08 = 256'h00000000000000000000000000000F0F0F0F0F0F0F0F00000000000000000000;
defparam rom_inst_0.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_0A = 256'h0000000000000000000000000000000000000F0F0F0F0F0F0F0F000000000000;
defparam rom_inst_0.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_0C = 256'h000000000000000000000000000000000000000000000F0F0F0F0F0F0F0F0000;
defparam rom_inst_0.INIT_RAM_0D = 256'h0F0F000000000000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_0E = 256'h00000000000000000000000000000000000000000000000000000F0F0F0F0F0F;
defparam rom_inst_0.INIT_RAM_0F = 256'h0F0F0F0F0F0F0000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000F0F;
defparam rom_inst_0.INIT_RAM_11 = 256'h00000F0F0F0F0F0F0F0F00000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_13 = 256'h0000000000000F0F0F0F0F0F0F0F000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_15 = 256'h000000000000000000000F0F0F0F0F0F0F0F0000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_17 = 256'h00000000000000000000000000000F0F0F0F0F0F0F0F00000000000000000000;
defparam rom_inst_0.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_19 = 256'h0000000000000000000000000000000000000F0F0F0F0F0F0F0F000000000000;
defparam rom_inst_0.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_1B = 256'h000000000000000000000000000000000000000000000F0F0F0F0F0F0F0F0000;
defparam rom_inst_0.INIT_RAM_1C = 256'h0F0F000000000000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_1D = 256'h00000000000000000000000000000000000000000000000000000F0F0F0F0F0F;
defparam rom_inst_0.INIT_RAM_1E = 256'h0F0F0F0F0F0F0000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000F0F;
defparam rom_inst_0.INIT_RAM_20 = 256'h00000F0F0F0F0F0F0F0F00000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_22 = 256'h0000000000000F0F0F0F0F0F0F0F000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_24 = 256'h000000000000000000000F0F0F0F0F0F0F0F0000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_26 = 256'h00000000000000000000000000000F0F0F0F0F0F0F0F00000000000000000000;
defparam rom_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000F0F0F0F0F0F0F0F000000000000;
defparam rom_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_2A = 256'h000000000000000000000000000000000000000000000F0F0F0F0F0F0F0F0000;
defparam rom_inst_0.INIT_RAM_2B = 256'h0F0F000000000000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_2C = 256'h00000000000000000000000000000000000000000000000000000F0F0F0F0F0F;
defparam rom_inst_0.INIT_RAM_2D = 256'h0F0F0F0F0F0F0000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000F0F;
defparam rom_inst_0.INIT_RAM_2F = 256'h00000F0F0F0F0F0F0F0F00000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_31 = 256'h0000000000000F0F0F0F0F0F0F0F000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_33 = 256'h000000000000000000000F0F0F0F0F0F0F0F0000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_35 = 256'h00000000000000000000000000000F0F0F0F0F0F0F0F00000000000000000000;
defparam rom_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam rom_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000F0F0F0F0F0F0F0F000000000000;
defparam rom_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //Gowin_ROM
